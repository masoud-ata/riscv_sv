typedef struct 
{
    logic [4:0] pc;
    logic [31:0] instruction;
} if_id_type;

